library verilog;
use verilog.vl_types.all;
entity testoperation is
end testoperation;
