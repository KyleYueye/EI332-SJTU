/////////////////////////////////////////////////////////////
//                                                         //
// School of Software of SJTU                              //
//                                                         //
/////////////////////////////////////////////////////////////

module sc_computer (resetn,mem_clk,pc,inst,aluout,memout,imem_clk,dmem_clk,in_port0,in_port1,out_port0,out_port1,out_port2,hex0,hex1,hex2,hex3,hex4,hex5);
   
   input resetn,mem_clk;
	reg clock;
	input [4:0] in_port0,in_port1;
   output [31:0] pc,inst,aluout,memout;
   output        imem_clk,dmem_clk;
	output [31:0] out_port0,out_port1,out_port2;
	output [6:0] hex0,hex1,hex2,hex3,hex4,hex5;
   wire   [31:0] data;
   wire          wmem; // all these "wire"s are used to connect or interface the cpu,dmem,imem and so on.
	
	always @(posedge mem_clk)
	begin
		if(~resetn)
			clock <= 0;
		clock <= ~clock;
	end
   
   sc_cpu cpu (clock,resetn,inst,memout,pc,wmem,aluout,data);          // CPU module.
   sc_instmem  imem (pc,inst,clock,mem_clk,imem_clk);                  // instruction memory.
   sc_datamem  dmem (aluout,data,memout,wmem,clock,mem_clk,dmem_clk,resetn,out_port0,out_port1,out_port2,in_port0,in_port1,mem_dataout,io_read_data); // data memory.

	sevenseg sevenseg0(out_port2[7:4],hex0);
	sevenseg sevenseg1(out_port2[3:0],hex1);
	sevenseg sevenseg2(out_port1[7:4],hex2);
	sevenseg sevenseg3(out_port1[3:0],hex3);
	sevenseg sevenseg4(out_port0[7:4],hex4);
	sevenseg sevenseg5(out_port0[3:0],hex5);

endmodule

module sevenseg ( data, ledsegments);
input [3:0] data;
output ledsegments;
reg [6:0] ledsegments;
always @ (*)
	case(data)
	// gfe_dcba // 7 段 LED 数码管的位段编号
	// 654_3210 // DE2 板上的信号位编号
		4'h0: ledsegments = 7'b100_0000; // DE2C 板上的数码管为共阳极接法。
		4'h1: ledsegments = 7'b111_1001;
		4'h2: ledsegments = 7'b010_0100;
		4'h3: ledsegments = 7'b011_0000;
		4'h4: ledsegments = 7'b001_1001;
		4'h5: ledsegments = 7'b001_0010;
		4'h6: ledsegments = 7'b000_0010;
		4'h7: ledsegments = 7'b111_1000;
		4'h8: ledsegments = 7'b000_0000;
		4'h9: ledsegments = 7'b001_0000;
		4'hA: ledsegments = 7'b000_1000;
		4'hB: ledsegments = 7'b000_0011;
		4'hC: ledsegments = 7'b100_0110;
		4'hD: ledsegments = 7'b010_0001;
		4'hE: ledsegments = 7'b000_0110;
		4'hF: ledsegments = 7'b000_1110;
		default: ledsegments = 7'b111_1111; // 其它值时全灭。
	endcase
endmodule



