library verilog;
use verilog.vl_types.all;
entity pipecomputer_sim is
end pipecomputer_sim;
